* HSPICE file created from 4NAND_f04.ext - technology: tsmc

.option scale=0.06u

M1000 Y1 Y Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=448 ps=208 
M1001 Vdd Y Y1 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 Y1 Y Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1003 Vdd Y Y1 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1004 a_9_68 Y gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=256 ps=104 
M1005 a_22_68 Y a_9_68 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1006 a_35_68 Y a_22_68 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1007 Y1 Y a_35_68 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1008 Y A Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=0 ps=0 
M1009 Vdd B Y Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1010 Y C Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1011 Vdd D Y Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1012 a_9_n30 A gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1013 a_22_n30 B a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1014 a_35_n30 C a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1015 Y D a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
C0 gnd Y 0.1fF
C1 gnd Y1 0.1fF
C2 Vdd Y 1.5fF
C3 Vdd Y1 0.6fF
C4 Y1 Y 0.0fF
C5 gnd gnd! 0.8fF
C6 Y1 gnd! 0.1fF
C7 Y gnd! 0.9fF
C8 Vdd gnd! 2.1fF

** hspice subcircuit dictionary
