magic
tech tsmc
timestamp 1492566096
<< nwell >>
rect -18 -8 39 16
<< ntransistor >>
rect 6 -22 9 -14
rect 19 -22 22 -14
<< ptransistor >>
rect 6 0 9 8
rect 19 0 22 8
<< ndiffusion >>
rect 0 -16 6 -14
rect 4 -22 6 -16
rect 9 -22 19 -14
rect 22 -22 75 -14
<< pdiffusion >>
rect 5 0 6 8
rect 9 0 10 8
rect 18 0 19 8
rect 22 0 23 8
<< ndcontact >>
rect -4 -24 4 -16
rect 75 -24 83 -16
<< pdcontact >>
rect -3 0 5 8
rect 10 0 18 8
rect 23 0 31 8
<< psubstratepcontact >>
rect 102 -32 110 -24
<< nsubstratencontact >>
rect -16 0 -8 8
<< polysilicon >>
rect 6 8 9 20
rect 19 8 22 20
rect 6 -14 9 0
rect 19 -14 22 0
rect 6 -26 9 -22
rect 19 -26 22 -22
<< polycontact >>
rect 4 20 12 28
rect 17 20 25 28
<< metal1 >>
rect -16 8 -12 43
rect -1 12 29 16
rect -1 8 3 12
rect 25 8 29 12
rect -8 0 -3 8
rect -16 -47 -12 0
rect 12 -4 16 0
rect 12 -8 81 -4
rect 77 -16 81 -8
rect 106 -24 110 43
rect -2 -28 2 -24
rect -2 -32 102 -28
rect 106 -47 110 -32
<< labels >>
rlabel metal1 -14 22 -14 22 3 Vdd
rlabel metal1 108 -9 108 -9 7 gnd
rlabel polysilicon 7 18 7 18 1 A
rlabel polysilicon 20 18 20 18 1 B
rlabel metal1 63 -6 63 -6 1 Y
<< end >>
