* SPICE3 file created from seg_a.ext - technology: tsmc

.option scale=0.06u
.include mosistsmc180.sp

V_paprika_0 D Gnd PULSE(0 3.3 2n 1n 1n 18n 40n)
V_paprika_1 C Gnd PULSE(0 3.3 2n 1n 1n 36n 80n)
V_paprika_2 B Gnd PULSE(0 3.3 2n 1n 1n 72n 160n)
V_paprika_3 A Gnd PULSE(0 3.3 2n 1n 1n 144n 320n)
V_paprika_4 Vdd Gnd DC 3.3

M1000 Y m1_24_n475 m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=152 pd=70 as=920 ps=422 
M1001 m1_0_86 m1_37_n478 Y m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 Y m1_49_n481 m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1003 x0/a_9_n26 m1_24_n475 m1_124_86 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=632 ps=286 
M1004 x0/a_22_n26 m1_37_n478 x0/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1005 Y m1_49_n481 x0/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1006 m1_49_n481 A m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1007 m1_0_86 B m1_49_n481 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1008 m1_49_n481 C m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1009 x1/a_9_n26 A m1_124_86 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1010 x1/a_22_n26 B x1/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1011 m1_49_n481 C x1/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1012 m1_37_n478 A m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1013 m1_0_86 B m1_37_n478 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1014 m1_37_n478 m1_35_n187 m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1015 x2/a_9_n26 A m1_124_86 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1016 x2/a_22_n26 B x2/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1017 m1_37_n478 m1_35_n187 x2/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1018 m1_24_n475 C m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=160 pd=72 as=0 ps=0 
M1019 m1_0_86 m1_35_n187 m1_24_n475 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1020 m1_24_n475 m1_48_n190 m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1021 m1_0_86 m1_66_n195 m1_24_n475 m1_0_86 pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1022 x3/a_9_n30 C m1_124_86 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1023 x3/a_22_n30 m1_35_n187 x3/a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1024 x3/a_35_n30 m1_48_n190 x3/a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1025 m1_24_n475 m1_66_n195 x3/a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1026 m1_35_n187 D m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1027 m1_35_n187 D m1_124_86 Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1028 m1_48_n190 B m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1029 m1_48_n190 B m1_124_86 Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1030 m1_66_n195 A m1_0_86 m1_0_86 pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1031 m1_66_n195 A m1_124_86 Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
C0 m1_48_n190 m1_24_n475 0.0fF
C1 m1_48_n190 m1_66_n195 4.5fF
C2 m1_24_n475 m1_49_n481 0.0fF
C3 m1_124_86 m1_37_n478 0.1fF
C4 m1_0_86 m1_35_n187 0.3fF
C5 m1_124_86 m1_48_n190 0.1fF
C6 m1_124_86 Y 0.1fF
C7 Y m1_37_n478 0.0fF
C8 m1_124_86 m1_49_n481 0.1fF
C9 m1_37_n478 m1_49_n481 0.5fF
C10 m1_0_86 m1_24_n475 0.8fF
C11 m1_0_86 m1_66_n195 0.3fF
C12 m1_24_n475 m1_35_n187 0.1fF
C13 Y m1_49_n481 0.0fF
C14 m1_35_n187 m1_66_n195 0.0fF
C15 m1_0_86 m1_37_n478 0.6fF
C16 m1_24_n475 m1_66_n195 0.0fF
C17 m1_124_86 m1_35_n187 0.1fF
C18 m1_37_n478 m1_35_n187 0.0fF
C19 m1_0_86 m1_48_n190 0.3fF
C20 Y m1_0_86 0.4fF
C21 m1_48_n190 m1_35_n187 4.8fF
C22 m1_0_86 m1_49_n481 0.5fF
C23 m1_124_86 m1_24_n475 0.1fF
C24 m1_24_n475 m1_37_n478 1.4fF
C25 m1_124_86 m1_66_n195 0.1fF
C26 m1_66_n195 GND 1.6fF
C27 m1_48_n190 GND 1.6fF
C28 m1_35_n187 GND 2.2fF
C29 m1_24_n475 GND 0.3fF
C30 m1_37_n478 GND 0.4fF
C31 m1_49_n481 GND 0.5fF
C32 m1_124_86 GND 2.6fF
C33 Y GND 0.1fF
C34 m1_0_86 GND 6.1fF

** hspice subcircuit dictionary
* x0	3NAND_2
* x1	3NAND_1
* x2	3NAND_0
* x3	4NAND_0

.tran 1n 320n

.control
set filetype=ascii
run
write segC.txt A B C D Y
.endc
.end
