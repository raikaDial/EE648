magic
tech tsmc
timestamp 1493235732
<< metal1 >>
rect -57 44 -53 86
rect -57 -560 -53 37
rect -46 -42 -42 86
rect -46 -368 -42 -49
rect -35 -128 -31 86
rect -46 -466 -42 -375
rect -35 -454 -31 -135
rect -24 -214 -20 86
rect 32 37 37 41
rect 148 40 152 86
rect 68 33 75 37
rect 31 -49 36 -45
rect 66 -53 75 -49
rect 31 -135 36 -131
rect 66 -139 75 -135
rect 31 -221 36 -217
rect -24 -274 -20 -221
rect 66 -225 75 -221
rect 37 -275 41 -269
rect 18 -281 22 -277
rect 55 -281 60 -277
rect -24 -442 -20 -281
rect 59 -313 75 -309
rect 37 -351 87 -347
rect 18 -375 24 -371
rect 37 -372 41 -351
rect 50 -363 87 -359
rect 50 -371 54 -363
rect 148 -368 152 33
rect 159 -46 163 86
rect 159 -274 163 -53
rect 170 -132 174 86
rect 170 -262 174 -139
rect 181 -218 185 86
rect 69 -375 87 -371
rect 72 -408 89 -404
rect -57 -740 -53 -567
rect -46 -740 -42 -473
rect -35 -548 -31 -461
rect -35 -740 -31 -555
rect -24 -740 -20 -449
rect 37 -466 41 -461
rect 49 -468 53 -449
rect 18 -473 24 -469
rect 60 -505 101 -501
rect 50 -555 111 -551
rect 37 -560 41 -555
rect 18 -566 22 -562
rect 50 -565 54 -555
rect 67 -567 111 -563
rect 73 -605 111 -601
rect 24 -633 75 -629
rect 24 -662 28 -633
rect 37 -644 87 -640
rect 37 -660 41 -644
rect 50 -653 99 -649
rect 50 -661 54 -653
rect 61 -663 111 -659
rect 148 -740 152 -375
rect 159 -560 163 -281
rect 170 -356 174 -269
rect 181 -344 185 -225
rect 159 -740 163 -567
rect 170 -740 174 -363
rect 181 -548 185 -351
rect 181 -740 185 -555
<< m2contact >>
rect -57 37 -50 44
rect -46 -49 -39 -42
rect -35 -135 -28 -128
rect -46 -375 -39 -368
rect 25 37 32 44
rect 75 33 82 40
rect 145 33 152 40
rect 24 -49 31 -42
rect 75 -53 82 -46
rect 24 -135 31 -128
rect 75 -139 82 -132
rect -24 -221 -17 -214
rect 24 -221 31 -214
rect 75 -225 82 -218
rect 36 -269 43 -262
rect -24 -281 -17 -274
rect 11 -281 18 -274
rect 60 -281 67 -274
rect 75 -316 82 -309
rect 87 -351 94 -344
rect 11 -375 18 -368
rect 87 -363 94 -356
rect 156 -53 163 -46
rect 167 -139 174 -132
rect 178 -225 185 -218
rect 167 -269 174 -262
rect 156 -281 163 -274
rect 87 -375 94 -368
rect 145 -375 152 -368
rect 89 -411 96 -404
rect -24 -449 -17 -442
rect 47 -449 54 -442
rect -35 -461 -28 -454
rect -46 -473 -39 -466
rect -57 -567 -50 -560
rect -35 -555 -28 -548
rect 35 -461 42 -454
rect 11 -473 18 -466
rect 101 -508 108 -501
rect 35 -555 42 -548
rect 111 -555 118 -548
rect 11 -567 18 -560
rect 111 -567 118 -560
rect 111 -608 118 -601
rect 75 -636 82 -629
rect 87 -644 94 -637
rect 99 -653 106 -646
rect 111 -663 118 -656
rect 178 -351 185 -344
rect 167 -363 174 -356
rect 158 -567 165 -560
rect 178 -555 185 -548
<< metal2 >>
rect -50 37 25 43
rect 82 33 145 38
rect -39 -49 24 -43
rect 82 -53 156 -48
rect -28 -135 24 -129
rect 82 -139 167 -134
rect -17 -221 24 -215
rect 82 -225 178 -220
rect 43 -269 167 -264
rect -17 -281 11 -276
rect 67 -281 156 -276
rect -39 -375 11 -370
rect -17 -449 47 -444
rect -28 -461 35 -456
rect -39 -473 11 -468
rect -28 -555 35 -550
rect -50 -567 11 -562
rect 77 -629 82 -316
rect 94 -351 178 -346
rect 94 -363 167 -358
rect 94 -375 145 -370
rect 89 -637 94 -411
rect 101 -646 106 -508
rect 118 -555 178 -550
rect 118 -567 158 -562
rect 113 -656 118 -608
use 1INV  1INV_0
timestamp 1493152604
transform 1 0 49 0 1 20
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493152604
transform 1 0 49 0 1 -66
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493152604
transform 1 0 49 0 1 -152
box -49 -20 79 66
use 1INV  1INV_3
timestamp 1493152604
transform 1 0 49 0 1 -238
box -49 -20 79 66
use 3NAND  3NAND_0
timestamp 1493160834
transform 1 0 18 0 1 -301
box -18 -51 110 43
use 4NAND  4NAND_0
timestamp 1493152043
transform 1 0 18 0 1 -395
box -18 -55 110 43
use 3NAND  3NAND_1
timestamp 1493160834
transform 1 0 18 0 1 -493
box -18 -51 110 43
use 4NAND  4NAND_1
timestamp 1493152043
transform 1 0 18 0 1 -587
box -18 -55 110 43
use 4NAND  4NAND_2
timestamp 1493152043
transform 1 0 18 0 1 -685
box -18 -55 110 43
<< labels >>
rlabel metal1 -57 -740 -53 86 3 A
rlabel metal1 -46 -740 -42 86 1 B
rlabel metal1 -35 -740 -31 86 1 C
rlabel metal1 -24 -740 -20 86 1 D
<< end >>
