magic
tech tsmc
timestamp 1492566197
<< nwell >>
rect -18 -8 52 16
<< ntransistor >>
rect 6 -26 9 -14
rect 19 -26 22 -14
rect 32 -26 35 -14
<< ptransistor >>
rect 6 0 9 8
rect 19 0 22 8
rect 32 0 35 8
<< ndiffusion >>
rect 0 -20 6 -14
rect 4 -26 6 -20
rect 9 -26 19 -14
rect 22 -26 32 -14
rect 35 -26 75 -14
<< pdiffusion >>
rect 5 0 6 8
rect 9 0 10 8
rect 18 0 19 8
rect 22 0 23 8
rect 31 0 32 8
rect 35 0 36 8
<< ndcontact >>
rect -4 -28 4 -20
rect 75 -28 83 -20
<< pdcontact >>
rect -3 0 5 8
rect 10 0 18 8
rect 23 0 31 8
rect 36 0 44 8
<< psubstratepcontact >>
rect 102 -36 110 -28
<< nsubstratencontact >>
rect -16 0 -8 8
<< polysilicon >>
rect 6 8 9 20
rect 19 8 22 20
rect 32 8 35 20
rect 6 -14 9 0
rect 19 -14 22 0
rect 32 -14 35 0
rect 6 -30 9 -26
rect 19 -30 22 -26
rect 32 -30 35 -26
<< polycontact >>
rect 4 20 12 28
rect 17 20 25 28
rect 30 20 38 28
<< metal1 >>
rect -16 8 -12 43
rect -1 12 29 16
rect -1 8 3 12
rect 25 8 29 12
rect -8 0 -3 8
rect -16 -51 -12 0
rect 12 -4 16 0
rect 38 -4 42 0
rect 12 -8 81 -4
rect 77 -20 81 -8
rect 106 -28 110 43
rect -2 -32 2 -28
rect -2 -36 102 -32
rect 106 -51 110 -36
<< labels >>
rlabel metal1 -14 22 -14 22 3 Vdd
rlabel metal1 108 -9 108 -9 7 gnd
rlabel polysilicon 7 18 7 18 1 A
rlabel polysilicon 20 18 20 18 1 B
rlabel polysilicon 33 18 33 18 1 C
rlabel metal1 68 -6 68 -6 1 Y
<< end >>
