magic
tech tsmc
timestamp 1492657465
<< nwell >>
rect -18 180 52 204
rect -18 86 52 110
rect -18 -8 52 16
<< ntransistor >>
rect 6 162 9 174
rect 19 162 22 174
rect 32 162 35 174
rect 6 68 9 80
rect 19 68 22 80
rect 32 68 35 80
rect 6 -26 9 -14
rect 19 -26 22 -14
rect 32 -26 35 -14
<< ptransistor >>
rect 6 188 9 196
rect 19 188 22 196
rect 32 188 35 196
rect 6 94 9 102
rect 19 94 22 102
rect 32 94 35 102
rect 6 0 9 8
rect 19 0 22 8
rect 32 0 35 8
<< ndiffusion >>
rect 0 170 6 174
rect 5 162 6 170
rect 9 162 19 174
rect 22 162 32 174
rect 35 170 44 174
rect 35 162 36 170
rect 0 76 6 80
rect 5 68 6 76
rect 9 68 19 80
rect 22 68 32 80
rect 35 76 44 80
rect 35 68 36 76
rect 0 -18 6 -14
rect 5 -26 6 -18
rect 9 -26 19 -14
rect 22 -26 32 -14
rect 35 -18 44 -14
rect 35 -26 36 -18
<< pdiffusion >>
rect 5 188 6 196
rect 9 188 10 196
rect 18 188 19 196
rect 22 188 23 196
rect 31 188 32 196
rect 35 188 36 196
rect 5 94 6 102
rect 9 94 10 102
rect 18 94 19 102
rect 22 94 23 102
rect 31 94 32 102
rect 35 94 36 102
rect 5 0 6 8
rect 9 0 10 8
rect 18 0 19 8
rect 22 0 23 8
rect 31 0 32 8
rect 35 0 36 8
<< ndcontact >>
rect -3 162 5 170
rect 36 162 44 170
rect -3 68 5 76
rect 36 68 44 76
rect -3 -26 5 -18
rect 36 -26 44 -18
<< pdcontact >>
rect -3 188 5 196
rect 10 188 18 196
rect 23 188 31 196
rect 36 188 44 196
rect -3 94 5 102
rect 10 94 18 102
rect 23 94 31 102
rect 36 94 44 102
rect -3 0 5 8
rect 10 0 18 8
rect 23 0 31 8
rect 36 0 44 8
<< psubstratepcontact >>
rect 102 152 110 160
rect 102 58 110 66
rect 102 -36 110 -28
<< nsubstratencontact >>
rect -16 188 -8 196
rect -16 94 -8 102
rect -16 0 -8 8
<< polysilicon >>
rect 6 196 9 208
rect 19 196 22 208
rect 32 196 35 208
rect 6 174 9 188
rect 19 174 22 188
rect 32 174 35 188
rect 6 158 9 162
rect 19 158 22 162
rect 32 158 35 162
rect 6 102 9 114
rect 19 102 22 114
rect 32 102 35 114
rect 6 80 9 94
rect 19 80 22 94
rect 32 80 35 94
rect 6 64 9 68
rect 19 64 22 68
rect 32 64 35 68
rect 6 8 9 20
rect 19 8 22 20
rect 32 8 35 20
rect 6 -14 9 0
rect 19 -14 22 0
rect 32 -14 35 0
rect 6 -30 9 -26
rect 19 -30 22 -26
rect 32 -30 35 -26
<< polycontact >>
rect 4 208 12 216
rect 17 208 25 216
rect 30 208 38 216
rect 4 114 12 122
rect 17 114 25 122
rect 30 114 38 122
rect 4 20 12 28
rect 17 20 25 28
rect 30 20 38 28
<< metal1 >>
rect -18 215 -14 231
rect -18 211 4 215
rect -18 196 -14 211
rect 25 211 30 215
rect 38 211 51 215
rect -1 200 29 204
rect -1 196 3 200
rect 25 196 29 200
rect -18 188 -16 196
rect -8 188 -3 196
rect -18 121 -14 188
rect 12 184 16 188
rect 38 184 42 188
rect 12 180 42 184
rect 38 170 42 180
rect -2 156 2 162
rect 106 160 110 231
rect -2 152 102 156
rect -18 117 4 121
rect -18 102 -14 117
rect 25 116 30 120
rect 38 116 50 120
rect -1 106 29 110
rect -1 102 3 106
rect 25 102 29 106
rect -18 94 -16 102
rect -8 94 -3 102
rect -18 8 -14 94
rect 12 90 16 94
rect 38 90 42 94
rect 12 86 42 90
rect 38 76 42 86
rect -2 62 2 68
rect 106 66 110 152
rect -2 58 102 62
rect 6 48 83 52
rect 6 28 10 48
rect 19 35 72 39
rect 19 28 23 35
rect 38 22 61 26
rect -1 12 29 16
rect -1 8 3 12
rect 25 8 29 12
rect -18 0 -16 8
rect -8 0 -3 8
rect -18 -51 -14 0
rect 12 -4 16 0
rect 38 -4 42 0
rect 12 -8 49 -4
rect 38 -18 42 -8
rect -2 -32 2 -26
rect 106 -28 110 58
rect -2 -36 102 -32
rect 106 -51 110 -36
rect 20 -119 24 -97
rect 50 -100 61 -96
rect 20 -123 32 -119
rect 19 -205 23 -183
rect 52 -187 72 -183
rect 19 -209 32 -205
rect 53 -274 83 -270
<< m2contact >>
rect 51 208 59 216
rect 50 113 58 121
rect 83 46 91 54
rect 72 33 80 41
rect 61 20 69 28
rect 49 -9 57 -1
rect 61 -102 69 -94
rect 72 -189 80 -181
rect 83 -276 91 -268
<< metal2 >>
rect 52 121 57 208
rect 51 -1 56 113
rect 63 -94 68 20
rect 74 -181 79 33
rect 85 -268 90 46
use 1INV  1INV_0
timestamp 1492656010
transform 1 0 31 0 1 -117
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1492656010
transform 1 0 31 0 1 -203
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1492656010
transform 1 0 31 0 1 -289
box -49 -20 79 66
<< labels >>
rlabel metal1 108 -9 108 -9 7 gnd
rlabel metal1 -16 22 -16 22 3 Vdd
rlabel metal1 108 85 108 85 7 gnd
rlabel metal1 -16 116 -16 116 3 Vdd
rlabel metal1 108 179 108 179 7 gnd
rlabel metal1 -16 210 -16 210 3 Vdd
rlabel metal1 12 86 42 90 1 Y1
rlabel metal1 12 180 42 184 1 Y2
rlabel space 18 -272 26 -264 1 stim
rlabel metal1 6 28 10 52 1 A
rlabel metal1 12 -8 49 -4 1 Y
<< end >>
