magic
tech tsmc
timestamp 1492568781
<< nwell >>
rect -18 -8 66 16
<< ntransistor >>
rect 6 -30 9 -14
rect 19 -30 22 -14
rect 32 -30 35 -14
rect 45 -30 48 -14
<< ptransistor >>
rect 6 0 9 8
rect 19 0 22 8
rect 32 0 35 8
rect 45 0 48 8
<< ndiffusion >>
rect 0 -22 6 -14
rect 4 -30 6 -22
rect 9 -30 19 -14
rect 22 -30 32 -14
rect 35 -30 45 -14
rect 48 -22 54 -14
rect 48 -30 49 -22
<< pdiffusion >>
rect 5 0 6 8
rect 9 0 10 8
rect 18 0 19 8
rect 22 0 23 8
rect 31 0 32 8
rect 35 0 36 8
rect 44 0 45 8
rect 48 0 49 8
<< ndcontact >>
rect -4 -30 4 -22
rect 49 -30 57 -22
<< pdcontact >>
rect -3 0 5 8
rect 10 0 18 8
rect 23 0 31 8
rect 36 0 44 8
rect 49 0 57 8
<< psubstratepcontact >>
rect 102 -40 110 -32
<< nsubstratencontact >>
rect -16 0 -8 8
<< polysilicon >>
rect 6 8 9 20
rect 19 8 22 20
rect 32 8 35 20
rect 45 8 48 20
rect 6 -14 9 0
rect 19 -14 22 0
rect 32 -14 35 0
rect 45 -14 48 0
rect 6 -34 9 -30
rect 19 -34 22 -30
rect 32 -34 35 -30
rect 45 -34 48 -30
<< polycontact >>
rect 4 20 12 28
rect 17 20 25 28
rect 30 20 38 28
rect 43 20 51 28
<< metal1 >>
rect -18 8 -14 43
rect -1 12 55 16
rect -1 8 3 12
rect 25 8 29 12
rect 51 8 55 12
rect -18 0 -16 8
rect -8 0 -3 8
rect -18 -55 -14 0
rect 12 -4 16 0
rect 38 -4 42 0
rect 12 -8 55 -4
rect 51 -22 55 -8
rect -2 -36 2 -30
rect 106 -32 110 43
rect -2 -40 102 -36
rect 106 -55 110 -40
<< labels >>
rlabel metal1 108 -9 108 -9 7 gnd
rlabel polysilicon 7 18 7 18 1 A
rlabel polysilicon 20 18 20 18 1 B
rlabel polysilicon 33 18 33 18 1 C
rlabel polysilicon 46 18 46 18 1 D
rlabel metal1 -16 22 -16 22 3 Vdd
rlabel metal1 52 -6 52 -6 1 Y
<< end >>
