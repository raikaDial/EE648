magic
tech tsmc
timestamp 1493154333
<< metal1 >>
rect -57 232 -53 531
rect -46 318 -42 531
rect -35 405 -31 531
rect -24 490 -20 531
rect 25 484 37 488
rect -57 -88 -53 225
rect -46 -12 -42 311
rect -57 -185 -53 -95
rect -57 -389 -53 -192
rect -46 -197 -42 -19
rect -35 -99 -31 398
rect -24 86 -20 483
rect 71 481 83 485
rect 24 398 36 402
rect 66 394 83 398
rect 24 312 36 316
rect 66 308 83 312
rect 24 226 36 230
rect 148 229 152 531
rect 159 315 163 531
rect 170 401 174 531
rect 181 488 185 531
rect 66 222 83 226
rect 18 80 23 84
rect 37 82 41 100
rect 50 84 54 90
rect 148 85 152 222
rect 159 97 163 308
rect 170 109 174 394
rect -46 -389 -42 -204
rect -35 -389 -31 -106
rect -24 -111 -20 79
rect 66 78 73 82
rect 73 42 77 46
rect 37 6 92 10
rect 18 -17 23 -13
rect 37 -14 41 6
rect 50 -6 92 -2
rect 50 -16 54 -6
rect 148 -14 152 78
rect 63 -18 92 -14
rect 73 -58 88 -54
rect 37 -110 41 -106
rect 50 -112 54 -95
rect 18 -116 23 -112
rect 69 -116 105 -112
rect -24 -209 -20 -118
rect 69 -155 100 -151
rect 18 -214 23 -210
rect 37 -215 41 -204
rect 50 -209 54 -193
rect 69 -214 112 -210
rect -24 -389 -20 -216
rect 69 -252 112 -248
rect 24 -282 75 -278
rect 24 -310 28 -282
rect 37 -294 87 -290
rect 37 -310 41 -294
rect 50 -302 100 -298
rect 50 -312 54 -302
rect 63 -312 112 -308
rect 148 -389 152 -21
rect 159 -110 163 90
rect 159 -389 163 -117
rect 170 -209 174 102
rect 181 11 185 481
rect 181 -2 185 4
rect 170 -389 174 -216
rect 181 -389 185 -9
<< m2contact >>
rect -24 483 -17 490
rect 18 483 25 490
rect -35 398 -28 405
rect -46 311 -39 318
rect -57 225 -50 232
rect -46 -19 -39 -12
rect -57 -95 -50 -88
rect -57 -192 -50 -185
rect 83 481 90 488
rect 17 397 24 404
rect 83 394 90 401
rect 17 311 24 318
rect 83 308 90 315
rect 17 225 24 232
rect 178 481 185 488
rect 167 394 174 401
rect 156 308 163 315
rect 83 222 90 229
rect 145 222 152 229
rect 36 100 43 107
rect -24 79 -17 86
rect 11 79 18 86
rect 49 90 56 97
rect 167 102 174 109
rect 156 90 163 97
rect -35 -106 -28 -99
rect -46 -204 -39 -197
rect 73 78 80 85
rect 145 78 152 85
rect 77 40 84 47
rect 11 -19 18 -12
rect 92 3 99 10
rect 92 -9 99 -2
rect 92 -21 99 -14
rect 145 -21 152 -14
rect 88 -61 95 -54
rect 49 -95 56 -88
rect 35 -106 42 -99
rect -24 -118 -17 -111
rect 11 -118 18 -111
rect 105 -117 112 -110
rect 100 -158 107 -151
rect 48 -193 55 -186
rect 35 -204 42 -197
rect -24 -216 -17 -209
rect 11 -216 18 -209
rect 112 -216 119 -209
rect 112 -255 119 -248
rect 75 -285 82 -278
rect 87 -294 94 -287
rect 100 -302 107 -295
rect 112 -313 119 -306
rect 156 -117 163 -110
rect 178 4 185 11
rect 178 -9 185 -2
rect 167 -216 174 -209
<< metal2 >>
rect -17 484 18 489
rect 90 482 178 487
rect -28 398 17 403
rect 90 395 167 400
rect -39 312 17 317
rect 90 309 156 314
rect -50 226 17 231
rect 90 223 145 228
rect 43 102 167 107
rect 56 91 156 96
rect -17 80 11 85
rect 80 79 145 84
rect -39 -18 11 -13
rect -50 -94 49 -89
rect -28 -105 35 -100
rect -17 -117 11 -112
rect -50 -192 48 -187
rect -39 -203 35 -198
rect -17 -215 11 -210
rect 77 -278 82 40
rect 99 4 178 9
rect 99 -8 178 -3
rect 99 -20 145 -15
rect 89 -287 94 -61
rect 112 -116 156 -111
rect 102 -295 107 -158
rect 119 -215 167 -210
rect 112 -306 117 -255
use 1INV  1INV_4
timestamp 1493152604
transform 1 0 49 0 1 465
box -49 -20 79 66
use 1INV  1INV_3
timestamp 1493152604
transform 1 0 49 0 1 379
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493152604
transform 1 0 49 0 1 293
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493152604
transform 1 0 49 0 1 207
box -49 -20 79 66
use 1INV  1INV_0
timestamp 1493152604
transform 1 0 49 0 1 121
box -49 -20 79 66
use 4NAND  4NAND_0
timestamp 1493152043
transform 1 0 18 0 1 58
box -18 -55 110 43
use 4NAND  4NAND_1
timestamp 1493152043
transform 1 0 18 0 1 -40
box -18 -55 110 43
use 4NAND  4NAND_2
timestamp 1493152043
transform 1 0 18 0 1 -138
box -18 -55 110 43
use 4NAND  4NAND_3
timestamp 1493152043
transform 1 0 18 0 1 -236
box -18 -55 110 43
use 4NAND  4NAND_4
timestamp 1493152043
transform 1 0 18 0 1 -334
box -18 -55 110 43
<< labels >>
rlabel metal1 -24 -389 -20 531 1 D
rlabel metal1 -35 -389 -31 531 1 C
rlabel metal1 -46 -389 -42 531 1 B
rlabel metal1 -57 -389 -53 531 3 A
<< end >>
