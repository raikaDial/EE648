magic
tech tsmc
timestamp 1493249081
<< metal1 >>
rect 0 86 4 93
rect 124 86 128 93
rect -57 44 -53 86
rect -57 -384 -53 37
rect -46 -188 -42 86
rect -35 -42 -31 86
rect -46 -290 -42 -195
rect -35 -278 -31 -49
rect -24 -128 -20 86
rect 148 41 152 86
rect 31 37 44 41
rect 66 34 75 38
rect 31 -49 44 -45
rect 66 -52 75 -48
rect 32 -135 44 -131
rect -24 -176 -20 -135
rect 66 -138 75 -134
rect -57 -480 -53 -391
rect -46 -468 -42 -297
rect -35 -372 -31 -285
rect -24 -360 -20 -183
rect 37 -187 41 -183
rect 49 -190 53 -183
rect 148 -188 152 34
rect 159 -45 163 86
rect 159 -176 163 -52
rect 170 -131 174 86
rect 18 -195 25 -191
rect 68 -195 73 -191
rect 69 -232 77 -228
rect 0 -275 4 -265
rect 124 -279 128 -266
rect 36 -289 40 -285
rect 18 -297 25 -293
rect 54 -297 87 -293
rect 58 -331 87 -327
rect -57 -658 -53 -487
rect -46 -658 -42 -475
rect -35 -658 -31 -379
rect -24 -658 -20 -367
rect 37 -383 41 -379
rect 50 -386 54 -367
rect 18 -391 23 -387
rect 56 -425 99 -421
rect 0 -466 4 -460
rect 124 -470 128 -459
rect 37 -481 41 -475
rect 18 -487 23 -483
rect 56 -487 111 -483
rect 56 -521 111 -517
rect 24 -553 77 -549
rect 0 -566 4 -557
rect 24 -578 28 -553
rect 37 -562 89 -558
rect 37 -579 41 -562
rect 124 -563 128 -554
rect 50 -570 101 -566
rect 50 -578 54 -570
rect 65 -581 111 -577
rect 69 -618 77 -614
rect 148 -658 152 -195
rect 159 -658 163 -183
rect 170 -290 174 -138
rect 170 -480 174 -297
rect 170 -658 174 -487
<< m2contact >>
rect -57 37 -50 44
rect -35 -49 -28 -42
rect -46 -195 -39 -188
rect 24 37 31 44
rect 75 34 82 41
rect 145 34 152 41
rect 24 -49 31 -42
rect 75 -52 82 -45
rect -24 -135 -17 -128
rect 25 -135 32 -128
rect 75 -138 82 -131
rect -24 -183 -17 -176
rect 35 -183 42 -176
rect 48 -183 55 -176
rect -35 -285 -28 -278
rect -46 -297 -39 -290
rect -57 -391 -50 -384
rect 11 -195 18 -188
rect 156 -52 163 -45
rect 167 -138 174 -131
rect 156 -183 163 -176
rect 73 -195 80 -188
rect 145 -195 152 -188
rect 77 -233 84 -226
rect 35 -285 42 -278
rect 11 -297 18 -290
rect 87 -297 94 -290
rect 87 -334 94 -327
rect -24 -367 -17 -360
rect 48 -367 55 -360
rect -35 -379 -28 -372
rect -46 -475 -39 -468
rect -57 -487 -50 -480
rect 35 -379 42 -372
rect 11 -391 18 -384
rect 99 -425 106 -418
rect 35 -475 42 -468
rect 11 -487 18 -480
rect 111 -487 118 -480
rect 111 -524 118 -517
rect 77 -554 84 -547
rect 89 -562 96 -555
rect 101 -570 108 -563
rect 111 -582 118 -575
rect 77 -621 84 -614
rect 167 -297 174 -290
rect 167 -487 174 -480
<< metal2 >>
rect -50 37 24 42
rect 82 34 145 39
rect -28 -49 24 -44
rect 82 -52 156 -47
rect -17 -135 25 -130
rect 82 -138 167 -133
rect -17 -183 35 -178
rect 55 -183 156 -178
rect -39 -195 11 -190
rect 80 -195 145 -190
rect -28 -285 35 -280
rect -39 -297 11 -292
rect -17 -367 48 -362
rect -28 -379 35 -374
rect -50 -391 11 -386
rect -39 -475 35 -470
rect -50 -487 11 -482
rect 77 -547 82 -233
rect 94 -297 167 -292
rect 89 -555 94 -334
rect 101 -563 106 -425
rect 118 -487 167 -482
rect 113 -575 118 -524
rect 79 -667 84 -621
use 1INV  1INV_0
timestamp 1493248008
transform 1 0 49 0 1 20
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493248008
transform 1 0 49 0 1 -66
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493248008
transform 1 0 49 0 1 -152
box -49 -20 79 66
use 4NAND  4NAND_0
timestamp 1493246152
transform 1 0 18 0 1 -215
box -18 -55 110 43
use 3NAND  3NAND_1
timestamp 1493246171
transform 1 0 18 0 1 -317
box -18 -51 110 43
use 3NAND  3NAND_0
timestamp 1493246171
transform 1 0 18 0 1 -411
box -18 -51 110 43
use 3NAND  3NAND_2
timestamp 1493246171
transform 1 0 18 0 1 -507
box -18 -51 110 43
use 4NAND  4NAND_3
timestamp 1493246152
transform 1 0 18 0 1 -603
box -18 -55 110 43
<< labels >>
rlabel metal1 -57 -658 -53 86 3 A
rlabel metal1 -46 -658 -42 86 1 B
rlabel metal1 -35 -658 -31 86 1 C
rlabel metal1 -24 -658 -20 86 1 D
rlabel metal1 0 86 4 93 5 Vdd
rlabel metal1 124 86 128 93 5 Gnd
rlabel metal2 79 -667 84 -662 1 Y
<< end >>
