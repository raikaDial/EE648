* HSPICE file created from seg_d.ext - technology: tsmc

.option scale=0.06u

M1000 Y m1_24_n662 Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=1296 ps=596 
M1001 Vdd m1_37_n660 Y Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 Y m1_50_n661 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1003 Vdd m1_61_n663 Y Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1004 x0/a_9_n30 m1_24_n662 Gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=864 ps=384 
M1005 x0/a_22_n30 m1_37_n660 x0/a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1006 x0/a_35_n30 m1_50_n661 x0/a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1007 Y m1_61_n663 x0/a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1008 m1_61_n663 A Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=0 ps=0 
M1009 Vdd C m1_61_n663 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1010 m1_61_n663 m1_37_n372 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1011 Vdd m1_55_n281 m1_61_n663 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1012 x1/a_9_n30 A Gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1013 x1/a_22_n30 C x1/a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1014 x1/a_35_n30 m1_37_n372 x1/a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1015 m1_61_n663 m1_55_n281 x1/a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1016 m1_50_n661 B Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1017 Vdd C m1_50_n661 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1018 m1_50_n661 D Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1019 x2/a_9_n26 B Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1020 x2/a_22_n26 C x2/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1021 m1_50_n661 D x2/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1022 m1_37_n660 B Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=0 ps=0 
M1023 Vdd m1_37_n372 m1_37_n660 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1024 m1_37_n660 m1_36_n269 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1025 Vdd m1_68_33 m1_37_n660 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1026 x3/a_9_n30 B Gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1027 x3/a_22_n30 m1_37_n372 x3/a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1028 x3/a_35_n30 m1_36_n269 x3/a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1029 m1_37_n660 m1_68_33 x3/a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1030 m1_24_n662 D Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1031 Vdd m1_36_n269 m1_24_n662 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1032 m1_24_n662 m1_55_n281 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1033 x4/a_9_n26 D Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1034 x4/a_22_n26 m1_36_n269 x4/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1035 m1_24_n662 m1_55_n281 x4/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1036 m1_37_n372 D Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1037 m1_37_n372 D Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1038 m1_36_n269 C Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1039 m1_36_n269 C Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1040 m1_55_n281 B Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1041 m1_55_n281 B Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1042 m1_68_33 A Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1043 m1_68_33 A Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
C0 m1_55_n281 Gnd 0.1fF
C1 m1_61_n663 m1_37_n372 0.0fF
C2 m1_50_n661 Vdd 0.6fF
C3 Y m1_50_n661 0.0fF
C4 m1_68_33 m1_37_n372 0.0fF
C5 m1_55_n281 m1_37_n372 0.6fF
C6 m1_36_n269 Gnd 0.1fF
C7 Y Gnd 0.1fF
C8 m1_61_n663 m1_55_n281 0.0fF
C9 m1_68_33 m1_55_n281 5.0fF
C10 m1_36_n269 m1_37_n372 5.8fF
C11 Vdd m1_37_n372 0.4fF
C12 m1_61_n663 Vdd 0.8fF
C13 m1_61_n663 Y 0.0fF
C14 m1_68_33 m1_36_n269 0.7fF
C15 m1_68_33 Vdd 0.3fF
C16 m1_36_n269 m1_55_n281 5.9fF
C17 m1_55_n281 Vdd 0.3fF
C18 m1_24_n662 m1_37_n660 2.0fF
C19 m1_36_n269 Vdd 0.4fF
C20 Y Vdd 0.6fF
C21 m1_37_n660 m1_50_n661 1.4fF
C22 m1_37_n660 Gnd 0.1fF
C23 m1_24_n662 m1_50_n661 0.0fF
C24 m1_37_n660 m1_37_n372 0.0fF
C25 m1_37_n660 m1_61_n663 0.0fF
C26 m1_24_n662 Gnd 0.1fF
C27 m1_68_33 m1_37_n660 0.0fF
C28 m1_37_n660 m1_55_n281 0.0fF
C29 m1_50_n661 Gnd 0.1fF
C30 m1_24_n662 m1_37_n372 0.1fF
C31 m1_24_n662 m1_61_n663 0.0fF
C32 m1_68_33 m1_24_n662 0.1fF
C33 m1_36_n269 m1_37_n660 0.0fF
C34 m1_37_n660 Vdd 0.8fF
C35 m1_37_n660 Y 0.0fF
C36 m1_50_n661 m1_37_n372 0.1fF
C37 m1_24_n662 m1_55_n281 0.0fF
C38 m1_61_n663 m1_50_n661 0.8fF
C39 Gnd m1_37_n372 0.1fF
C40 m1_61_n663 Gnd 0.1fF
C41 m1_55_n281 m1_50_n661 0.1fF
C42 m1_24_n662 m1_36_n269 0.1fF
C43 m1_24_n662 Vdd 0.6fF
C44 m1_68_33 Gnd 0.1fF
C45 m1_68_33 gnd! 2.0fF
C46 m1_55_n281 gnd! 2.3fF
C47 m1_36_n269 gnd! 2.4fF
C48 m1_37_n372 gnd! 2.7fF
C49 m1_24_n662 gnd! 0.3fF
C50 m1_37_n660 gnd! 0.3fF
C51 m1_50_n661 gnd! 0.5fF
C52 m1_61_n663 gnd! 0.5fF
C53 Gnd gnd! 3.4fF
C54 Y gnd! 0.1fF
C55 Vdd gnd! 7.9fF

** hspice subcircuit dictionary
* x0	4NAND_2
* x1	4NAND_1
* x2	3NAND_1
* x3	4NAND_0
* x4	3NAND_0
