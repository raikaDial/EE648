magic
tech tsmc
timestamp 1493254982
<< metal1 >>
rect 0 87 4 97
rect 124 87 128 97
rect -57 45 -53 87
rect -57 -445 -53 38
rect -46 -41 -42 87
rect -57 -552 -53 -452
rect -46 -457 -42 -48
rect -35 -127 -31 87
rect -35 -280 -31 -134
rect -24 -187 -20 87
rect 148 44 152 89
rect 32 38 38 42
rect 70 38 75 43
rect 32 -48 39 -44
rect 69 -48 75 -43
rect 32 -134 41 -130
rect 68 -135 75 -130
rect 148 -174 152 37
rect 159 -42 163 89
rect 37 -188 41 -182
rect 18 -194 26 -189
rect 54 -194 60 -189
rect -35 -360 -31 -287
rect -46 -552 -42 -464
rect -35 -552 -31 -367
rect -24 -375 -20 -194
rect 56 -226 75 -222
rect 148 -267 152 -181
rect 159 -187 163 -49
rect 170 -128 174 89
rect 37 -274 90 -269
rect 37 -284 42 -274
rect 18 -288 25 -284
rect 54 -286 90 -281
rect 59 -320 87 -314
rect 37 -377 42 -368
rect 148 -375 152 -274
rect 159 -279 163 -194
rect 18 -381 24 -377
rect 54 -382 99 -377
rect -24 -469 -20 -382
rect 59 -414 101 -410
rect 37 -470 41 -464
rect 50 -470 54 -452
rect 69 -464 113 -459
rect 63 -470 68 -464
rect 18 -475 24 -471
rect -24 -552 -20 -476
rect 69 -512 112 -508
rect 24 -542 76 -538
rect 24 -571 28 -542
rect 37 -554 88 -550
rect 148 -550 152 -382
rect 159 -550 163 -286
rect 170 -457 174 -135
rect 170 -550 174 -464
rect 37 -570 42 -554
rect 50 -562 100 -558
rect 50 -568 54 -562
rect 67 -573 112 -569
rect 71 -610 77 -606
<< m2contact >>
rect -57 38 -50 45
rect -46 -48 -39 -41
rect -57 -452 -50 -445
rect -35 -134 -28 -127
rect 25 38 32 45
rect 75 37 82 44
rect 145 37 152 44
rect 25 -48 32 -41
rect 75 -49 82 -42
rect 25 -134 32 -127
rect 75 -135 82 -128
rect 157 -49 164 -42
rect 36 -182 43 -175
rect 145 -181 152 -174
rect -24 -194 -17 -187
rect 11 -194 18 -187
rect 60 -194 67 -187
rect -35 -287 -28 -280
rect -35 -367 -28 -360
rect -46 -464 -39 -457
rect 75 -226 82 -219
rect 169 -135 176 -128
rect 156 -194 163 -187
rect 90 -274 97 -267
rect 145 -274 152 -267
rect 11 -288 18 -281
rect 90 -286 97 -279
rect 87 -320 94 -313
rect 36 -368 43 -361
rect -24 -382 -17 -375
rect 11 -382 18 -375
rect 156 -286 163 -279
rect 99 -382 106 -375
rect 145 -382 152 -375
rect 101 -415 108 -408
rect 48 -452 55 -445
rect 35 -464 42 -457
rect -24 -476 -17 -469
rect 11 -476 18 -469
rect 62 -464 69 -457
rect 113 -464 120 -457
rect 112 -513 119 -506
rect 76 -545 83 -538
rect 88 -554 95 -547
rect 167 -464 174 -457
rect 100 -562 107 -555
rect 112 -573 119 -566
rect 77 -612 84 -605
<< metal2 >>
rect -50 38 25 43
rect 82 37 145 42
rect -39 -48 25 -43
rect 82 -49 157 -44
rect -28 -134 25 -129
rect 82 -135 169 -130
rect 43 -181 145 -176
rect -17 -194 11 -189
rect 67 -194 156 -189
rect -28 -287 11 -282
rect -28 -367 36 -362
rect -17 -382 11 -377
rect -50 -452 48 -447
rect -39 -464 35 -459
rect -17 -475 11 -470
rect 77 -538 82 -226
rect 97 -274 145 -269
rect 97 -286 156 -281
rect 89 -547 94 -320
rect 106 -382 145 -377
rect 101 -555 106 -415
rect 120 -464 167 -459
rect 112 -566 117 -513
rect 79 -655 84 -612
use 1INV  1INV_0
timestamp 1493248008
transform 1 0 49 0 1 21
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493248008
transform 1 0 49 0 1 -65
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493248008
transform 1 0 49 0 1 -151
box -49 -20 79 66
use 3NAND  3NAND_0
timestamp 1493246171
transform 1 0 18 0 1 -214
box -18 -51 110 43
use 3NAND  3NAND_1
timestamp 1493246171
transform 1 0 18 0 1 -308
box -18 -51 110 43
use 3NAND  3NAND_2
timestamp 1493246171
transform 1 0 18 0 1 -402
box -18 -51 110 43
use 4NAND  4NAND_0
timestamp 1493246152
transform 1 0 18 0 1 -496
box -18 -55 110 43
use 4NAND  4NAND_1
timestamp 1493246152
transform 1 0 18 0 1 -594
box -18 -55 110 43
<< labels >>
rlabel metal1 -24 77 -20 87 1 D
rlabel metal1 -35 77 -31 87 1 C
rlabel metal1 -46 77 -42 87 1 B
rlabel metal1 -57 77 -53 87 3 A
rlabel metal1 0 87 4 97 5 Vdd
rlabel metal1 124 87 128 97 5 Gnd
rlabel metal2 79 -655 84 -650 1 Y
<< end >>
