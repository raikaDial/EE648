magic
tech tsmc
timestamp 1492568499
<< nwell >>
rect -16 -8 41 16
<< ntransistor >>
rect 8 -22 11 -14
rect 21 -22 24 -14
<< ptransistor >>
rect 8 0 11 8
rect 21 0 24 8
<< ndiffusion >>
rect 7 -22 8 -14
rect 11 -22 21 -14
rect 24 -22 25 -14
<< pdiffusion >>
rect 7 0 8 8
rect 11 0 12 8
rect 20 0 21 8
rect 24 0 25 8
<< ndcontact >>
rect -1 -22 7 -14
rect 25 -22 33 -14
<< pdcontact >>
rect -1 0 7 8
rect 12 0 20 8
rect 25 0 33 8
<< psubstratepcontact >>
rect 104 -32 112 -24
<< nsubstratencontact >>
rect -14 0 -6 8
<< polysilicon >>
rect 8 8 11 20
rect 21 8 24 20
rect 8 -14 11 0
rect 21 -14 24 0
rect 8 -26 11 -22
rect 21 -26 24 -22
<< polycontact >>
rect 6 20 14 28
rect 19 20 27 28
<< metal1 >>
rect -16 8 -12 43
rect 1 12 31 16
rect 1 8 5 12
rect 27 8 31 12
rect -16 0 -14 8
rect -6 0 -1 8
rect -16 -47 -12 0
rect 14 -4 18 0
rect 14 -8 31 -4
rect 27 -14 31 -8
rect 0 -28 4 -22
rect 108 -24 112 43
rect 0 -32 104 -28
rect 108 -47 112 -32
<< labels >>
rlabel polysilicon 9 18 9 18 1 A
rlabel polysilicon 22 18 22 18 1 B
rlabel metal1 -14 22 -14 22 3 Vdd
rlabel metal1 110 -9 110 -9 7 gnd
rlabel metal1 29 -10 29 -10 1 Y
<< end >>
