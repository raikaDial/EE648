magic
tech tsmc
timestamp 1493412550
<< metal1 >>
rect 57 843 61 869
rect 181 842 185 858
rect 319 845 323 869
rect 443 843 447 858
rect 570 844 574 869
rect 694 844 698 858
rect 821 844 825 869
rect 945 844 949 858
rect 1083 844 1087 869
rect 1207 844 1211 858
rect 1334 846 1338 869
rect 1458 846 1462 858
rect 1584 845 1588 869
rect 1708 844 1712 858
rect 1139 246 1153 250
rect 630 239 640 243
rect 388 131 398 135
rect 130 46 136 50
rect 0 -11 4 8
rect 11 -24 15 7
rect 22 -37 26 7
rect 33 -50 37 8
rect 136 -70 140 8
rect 262 -11 266 94
rect 273 -24 277 94
rect 284 -37 288 95
rect 295 -50 299 95
rect 398 -71 402 93
rect 513 -11 517 200
rect 524 -24 528 201
rect 535 -37 539 200
rect 546 -50 550 203
rect 640 -70 644 201
rect 894 50 908 54
rect 764 -11 768 12
rect 775 -24 779 12
rect 786 -37 790 13
rect 797 -50 801 13
rect 908 -70 912 12
rect 1026 -11 1030 208
rect 1037 -24 1041 208
rect 1048 -37 1052 208
rect 1059 -50 1063 208
rect 1153 -70 1157 208
rect 1277 -11 1281 200
rect 1288 -24 1292 199
rect 1299 -37 1303 200
rect 1310 -50 1314 201
rect 1403 139 1417 143
rect 1417 -70 1421 101
rect 1527 -11 1531 265
rect 1538 -24 1542 264
rect 1549 -37 1553 264
rect 1560 -50 1564 265
rect 1640 150 1654 154
rect 1654 -70 1658 112
<< m2contact >>
rect 57 869 64 876
rect 319 869 326 876
rect 570 869 577 876
rect 821 869 828 876
rect 1083 869 1090 876
rect 1334 869 1341 876
rect 1584 869 1591 876
rect 181 858 188 865
rect 443 858 450 865
rect 694 858 701 865
rect 945 858 952 865
rect 1207 858 1214 865
rect 1458 858 1465 865
rect 1708 858 1715 865
rect 1153 243 1160 250
rect 640 236 647 243
rect 1153 208 1160 215
rect 398 128 405 135
rect 136 43 143 50
rect 136 8 143 15
rect 0 -18 7 -11
rect 11 -31 18 -24
rect 22 -44 29 -37
rect 33 -57 40 -50
rect 262 -18 269 -11
rect 273 -31 280 -24
rect 284 -44 291 -37
rect 398 93 405 100
rect 295 -57 302 -50
rect 513 -18 520 -11
rect 524 -31 531 -24
rect 535 -44 542 -37
rect 640 201 647 208
rect 546 -57 553 -50
rect 908 47 915 54
rect 764 -18 771 -11
rect 775 -31 782 -24
rect 786 -44 793 -37
rect 908 12 915 19
rect 797 -57 804 -50
rect 1026 -18 1033 -11
rect 1037 -31 1044 -24
rect 1048 -44 1055 -37
rect 1059 -57 1066 -50
rect 1277 -18 1284 -11
rect 1288 -31 1295 -24
rect 1299 -44 1306 -37
rect 1417 136 1424 143
rect 1417 101 1424 108
rect 1310 -57 1317 -50
rect 1527 -18 1534 -11
rect 1538 -31 1545 -24
rect 1549 -44 1556 -37
rect 1654 147 1661 154
rect 1654 112 1661 119
rect 1560 -57 1567 -50
<< metal2 >>
rect 0 871 57 876
rect 64 871 319 876
rect 326 871 570 876
rect 577 871 821 876
rect 828 871 1083 876
rect 1090 871 1334 876
rect 1341 871 1584 876
rect 1591 871 1769 876
rect 0 858 181 863
rect 188 858 443 863
rect 450 858 694 863
rect 701 858 945 863
rect 952 858 1207 863
rect 1214 858 1458 863
rect 1465 858 1708 863
rect 1715 858 1769 863
rect 640 208 646 236
rect 1153 215 1159 243
rect 398 100 404 128
rect 1417 108 1423 136
rect 1654 119 1660 147
rect 136 15 142 43
rect 908 19 914 47
rect 7 -18 262 -13
rect 269 -18 513 -13
rect 520 -18 764 -13
rect 771 -18 1026 -13
rect 1033 -18 1277 -13
rect 1284 -18 1527 -13
rect 1534 -18 1769 -13
rect 0 -31 11 -26
rect 18 -31 273 -26
rect 280 -31 524 -26
rect 531 -31 775 -26
rect 782 -31 1037 -26
rect 1044 -31 1288 -26
rect 1295 -31 1538 -26
rect 1545 -31 1769 -26
rect 0 -44 22 -39
rect 29 -44 284 -39
rect 291 -44 535 -39
rect 542 -44 786 -39
rect 793 -44 1048 -39
rect 1055 -44 1299 -39
rect 1306 -44 1549 -39
rect 1556 -44 1769 -39
rect 0 -57 33 -52
rect 40 -57 295 -52
rect 302 -57 546 -52
rect 553 -57 797 -52
rect 804 -57 1059 -52
rect 1066 -57 1310 -52
rect 1317 -57 1560 -52
rect 1567 -57 1769 -52
use seg_a  seg_a_0
timestamp 1493411817
transform 1 0 57 0 1 307
box -57 -300 185 536
use seg_b  seg_b_0
timestamp 1493411841
transform 1 0 319 0 1 752
box -57 -658 174 93
use seg_c  seg_c_0
timestamp 1493411856
transform 1 0 570 0 1 752
box -57 -552 174 92
use seg_d  seg_d_0
timestamp 1493411876
transform 1 0 821 0 1 752
box -57 -740 185 92
use seg_e  seg_e_0
timestamp 1493411891
transform 1 0 1083 0 1 752
box -57 -544 174 92
use seg_f  seg_f_0
timestamp 1493411906
transform 1 0 1334 0 1 751
box -57 -649 176 97
use seg_g  seg_g_0
timestamp 1493411924
transform 1 0 1584 0 1 754
box -57 -642 185 93
<< labels >>
rlabel metal1 136 -70 140 8 1 seg_a
rlabel metal1 398 -71 402 93 1 seg_b
rlabel metal1 640 -70 644 201 1 seg_c
rlabel metal1 908 -70 912 12 1 seg_d
rlabel metal1 1153 -70 1157 208 1 seg_e
rlabel metal1 1417 -70 1421 101 1 seg_f
rlabel metal1 1654 -70 1658 112 1 seg_g
rlabel metal2 7 -18 262 -13 1 A
rlabel metal2 18 -31 273 -26 1 B
rlabel metal2 29 -44 284 -39 1 C
rlabel metal2 40 -57 295 -52 1 D
rlabel metal2 0 871 57 876 5 Vdd
rlabel metal2 0 858 181 863 1 Gnd
<< end >>
