magic
tech tsmc
timestamp 1493247679
<< metal1 >>
rect 0 531 4 536
rect 124 531 128 536
rect -57 232 -53 531
rect -46 318 -42 531
rect -35 405 -31 531
rect -24 490 -20 531
rect 25 484 37 488
rect -57 1 -53 225
rect -46 77 -42 311
rect -57 -96 -53 -6
rect -57 -300 -53 -103
rect -46 -108 -42 70
rect -35 -10 -31 398
rect -24 175 -20 483
rect 67 481 83 485
rect 24 398 36 402
rect 66 394 83 398
rect 24 312 36 316
rect 66 308 83 312
rect 24 226 36 230
rect 148 229 152 531
rect 159 315 163 531
rect 170 401 174 531
rect 181 488 185 531
rect 66 222 83 226
rect 18 169 23 173
rect 37 171 41 189
rect 50 173 54 179
rect 148 174 152 222
rect 159 186 163 308
rect 170 198 174 394
rect -46 -300 -42 -115
rect -35 -300 -31 -17
rect -24 -22 -20 168
rect 66 167 73 171
rect 73 131 77 135
rect 37 95 92 99
rect 18 72 23 76
rect 37 75 41 95
rect 50 83 92 87
rect 50 73 54 83
rect 148 75 152 167
rect 63 71 92 75
rect 73 31 88 35
rect 37 -21 41 -17
rect 50 -23 54 -6
rect 18 -27 23 -23
rect 69 -27 105 -23
rect -24 -120 -20 -29
rect 69 -66 100 -62
rect 18 -125 23 -121
rect 37 -126 41 -115
rect 50 -120 54 -104
rect 69 -125 112 -121
rect -24 -300 -20 -127
rect 69 -163 112 -159
rect 24 -193 75 -189
rect 24 -221 28 -193
rect 37 -205 87 -201
rect 37 -221 41 -205
rect 50 -213 100 -209
rect 50 -223 54 -213
rect 63 -223 112 -219
rect 148 -300 152 68
rect 159 -21 163 179
rect 159 -300 163 -28
rect 170 -120 174 191
rect 181 100 185 481
rect 181 87 185 93
rect 170 -300 174 -127
rect 181 -300 185 80
<< m2contact >>
rect -24 483 -17 490
rect 18 483 25 490
rect -35 398 -28 405
rect -46 311 -39 318
rect -57 225 -50 232
rect -46 70 -39 77
rect -57 -6 -50 1
rect -57 -103 -50 -96
rect 83 481 90 488
rect 17 397 24 404
rect 83 394 90 401
rect 17 311 24 318
rect 83 308 90 315
rect 17 225 24 232
rect 178 481 185 488
rect 167 394 174 401
rect 156 308 163 315
rect 83 222 90 229
rect 145 222 152 229
rect 36 189 43 196
rect -24 168 -17 175
rect 11 168 18 175
rect 49 179 56 186
rect 167 191 174 198
rect 156 179 163 186
rect -35 -17 -28 -10
rect -46 -115 -39 -108
rect 73 167 80 174
rect 145 167 152 174
rect 77 129 84 136
rect 11 70 18 77
rect 92 92 99 99
rect 92 80 99 87
rect 92 68 99 75
rect 145 68 152 75
rect 88 28 95 35
rect 49 -6 56 1
rect 35 -17 42 -10
rect -24 -29 -17 -22
rect 11 -29 18 -22
rect 105 -28 112 -21
rect 100 -69 107 -62
rect 48 -104 55 -97
rect 35 -115 42 -108
rect -24 -127 -17 -120
rect 11 -127 18 -120
rect 112 -127 119 -120
rect 112 -166 119 -159
rect 75 -196 82 -189
rect 87 -205 94 -198
rect 100 -213 107 -206
rect 112 -224 119 -217
rect 156 -28 163 -21
rect 178 93 185 100
rect 178 80 185 87
rect 167 -127 174 -120
<< metal2 >>
rect -17 484 18 489
rect 90 482 178 487
rect -28 398 17 403
rect 90 395 167 400
rect -39 312 17 317
rect 90 309 156 314
rect -50 226 17 231
rect 90 223 145 228
rect 43 191 167 196
rect 56 180 156 185
rect -17 169 11 174
rect 80 168 145 173
rect -39 71 11 76
rect -50 -5 49 0
rect -28 -16 35 -11
rect -17 -28 11 -23
rect -50 -103 48 -98
rect -39 -114 35 -109
rect -17 -126 11 -121
rect 77 -189 82 129
rect 99 93 178 98
rect 99 81 178 86
rect 99 69 145 74
rect 89 -198 94 28
rect 112 -27 156 -22
rect 102 -206 107 -69
rect 119 -126 167 -121
rect 112 -217 117 -166
use 1INV  1INV_4
timestamp 1493247659
transform 1 0 49 0 1 465
box -49 -20 79 66
use 1INV  1INV_3
timestamp 1493247659
transform 1 0 49 0 1 379
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493247659
transform 1 0 49 0 1 293
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493247659
transform 1 0 49 0 1 207
box -49 -20 79 66
use 4NAND  4NAND_0
timestamp 1493246152
transform 1 0 18 0 1 145
box -18 -55 110 43
use 4NAND  4NAND_1
timestamp 1493246152
transform 1 0 18 0 1 48
box -18 -55 110 43
use 4NAND  4NAND_2
timestamp 1493246152
transform 1 0 18 0 1 -49
box -18 -55 110 43
use 4NAND  4NAND_3
timestamp 1493246152
transform 1 0 18 0 1 -147
box -18 -55 110 43
use 4NAND  4NAND_4
timestamp 1493246152
transform 1 0 18 0 1 -245
box -18 -55 110 43
<< labels >>
rlabel metal1 -57 526 -53 531 4 A
rlabel metal1 -46 526 -42 531 5 B
rlabel metal1 -35 526 -31 531 5 C
rlabel metal1 -24 526 -20 531 5 D
rlabel metal1 0 531 4 536 5 Vdd
rlabel metal1 124 531 128 536 5 Gnd
<< end >>
