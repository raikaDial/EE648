magic
tech tsmc
timestamp 1492639596
<< nwell >>
rect -18 90 66 114
rect -18 -8 66 16
<< ntransistor >>
rect 6 68 9 84
rect 19 68 22 84
rect 32 68 35 84
rect 45 68 48 84
rect 6 -30 9 -14
rect 19 -30 22 -14
rect 32 -30 35 -14
rect 45 -30 48 -14
<< ptransistor >>
rect 6 98 9 106
rect 19 98 22 106
rect 32 98 35 106
rect 45 98 48 106
rect 6 0 9 8
rect 19 0 22 8
rect 32 0 35 8
rect 45 0 48 8
<< ndiffusion >>
rect 0 76 6 84
rect 4 68 6 76
rect 9 68 19 84
rect 22 68 32 84
rect 35 68 45 84
rect 48 76 54 84
rect 48 68 49 76
rect 0 -22 6 -14
rect 4 -30 6 -22
rect 9 -30 19 -14
rect 22 -30 32 -14
rect 35 -30 45 -14
rect 48 -22 54 -14
rect 48 -30 49 -22
<< pdiffusion >>
rect 5 98 6 106
rect 9 98 10 106
rect 18 98 19 106
rect 22 98 23 106
rect 31 98 32 106
rect 35 98 36 106
rect 44 98 45 106
rect 48 98 49 106
rect 5 0 6 8
rect 9 0 10 8
rect 18 0 19 8
rect 22 0 23 8
rect 31 0 32 8
rect 35 0 36 8
rect 44 0 45 8
rect 48 0 49 8
<< ndcontact >>
rect -4 68 4 76
rect 49 68 57 76
rect -4 -30 4 -22
rect 49 -30 57 -22
<< pdcontact >>
rect -3 98 5 106
rect 10 98 18 106
rect 23 98 31 106
rect 36 98 44 106
rect 49 98 57 106
rect -3 0 5 8
rect 10 0 18 8
rect 23 0 31 8
rect 36 0 44 8
rect 49 0 57 8
<< psubstratepcontact >>
rect 102 58 110 66
rect 102 -40 110 -32
<< nsubstratencontact >>
rect -16 98 -8 106
rect -16 0 -8 8
<< polysilicon >>
rect 6 106 9 118
rect 19 106 22 118
rect 32 106 35 118
rect 45 106 48 118
rect 6 84 9 98
rect 19 84 22 98
rect 32 84 35 98
rect 45 84 48 98
rect 6 64 9 68
rect 19 64 22 68
rect 32 64 35 68
rect 45 64 48 68
rect 6 8 9 20
rect 19 8 22 20
rect 32 8 35 20
rect 45 8 48 20
rect 6 -14 9 0
rect 19 -14 22 0
rect 32 -14 35 0
rect 45 -14 48 0
rect 6 -34 9 -30
rect 19 -34 22 -30
rect 32 -34 35 -30
rect 45 -34 48 -30
<< polycontact >>
rect 4 118 12 126
rect 17 118 25 126
rect 30 118 38 126
rect 43 118 51 126
rect 4 20 12 28
rect 17 20 25 28
rect 30 20 38 28
rect 43 20 51 28
<< metal1 >>
rect -18 106 -14 141
rect 12 120 17 124
rect 25 120 30 124
rect 38 120 43 124
rect 51 120 75 124
rect -1 110 55 114
rect -1 106 3 110
rect 25 106 29 110
rect 51 106 55 110
rect -18 98 -16 106
rect -8 98 -3 106
rect -18 8 -14 98
rect 12 94 16 98
rect 38 94 42 98
rect 12 90 55 94
rect 51 76 55 90
rect -2 62 2 68
rect 106 66 110 141
rect -2 58 102 62
rect -1 12 55 16
rect -1 8 3 12
rect 25 8 29 12
rect 51 8 55 12
rect -18 0 -16 8
rect -8 0 -3 8
rect -18 -55 -14 0
rect 12 -4 16 0
rect 38 -4 42 0
rect 12 -8 75 -4
rect 51 -22 55 -8
rect -2 -36 2 -30
rect 106 -32 110 58
rect -2 -40 102 -36
rect 106 -55 110 -40
<< m2contact >>
rect 75 117 83 125
rect 75 -10 83 -2
<< metal2 >>
rect 77 -2 82 117
<< labels >>
rlabel metal1 108 -9 108 -9 7 gnd
rlabel polysilicon 7 18 7 18 1 A
rlabel polysilicon 20 18 20 18 1 B
rlabel polysilicon 33 18 33 18 1 C
rlabel polysilicon 46 18 46 18 1 D
rlabel metal1 -16 22 -16 22 3 Vdd
rlabel metal1 52 -6 52 -6 1 Y
rlabel metal1 108 89 108 89 7 gnd
rlabel metal1 -16 120 -16 120 3 Vdd
rlabel metal1 51 76 55 94 1 Y1
<< end >>
