magic
tech tsmc
timestamp 1493192020
<< metal1 >>
rect -57 44 -53 86
rect -57 -286 -53 37
rect -46 -42 -42 86
rect -46 -274 -42 -49
rect -35 -188 -31 86
rect -24 -128 -20 86
rect 32 37 36 41
rect 148 40 152 86
rect 71 33 75 37
rect 32 -49 36 -45
rect 66 -53 75 -49
rect 32 -135 36 -131
rect -57 -380 -53 -293
rect -46 -368 -42 -281
rect -35 -356 -31 -195
rect -57 -552 -53 -387
rect -46 -552 -42 -375
rect -35 -552 -31 -363
rect -24 -552 -20 -135
rect 66 -139 75 -135
rect 35 -187 39 -173
rect 48 -190 52 -183
rect 148 -188 152 33
rect 159 -46 163 86
rect 159 -176 163 -53
rect 170 -132 174 86
rect 170 -164 174 -139
rect 18 -195 23 -191
rect 66 -195 73 -191
rect 72 -233 77 -229
rect 37 -286 41 -281
rect 18 -293 24 -289
rect 52 -293 89 -289
rect 59 -326 89 -322
rect 18 -386 27 -382
rect 36 -386 40 -375
rect 50 -379 54 -365
rect 60 -419 101 -415
rect 24 -451 77 -447
rect 24 -475 28 -451
rect 37 -462 89 -458
rect 37 -478 41 -462
rect 49 -481 101 -477
rect 148 -552 152 -195
rect 159 -552 163 -183
rect 170 -286 174 -171
rect 170 -552 174 -293
<< m2contact >>
rect -57 37 -50 44
rect -46 -49 -39 -42
rect 25 37 32 44
rect 75 33 82 40
rect 145 33 152 40
rect 25 -49 32 -42
rect 75 -53 82 -46
rect -24 -135 -17 -128
rect 25 -135 32 -128
rect -35 -195 -28 -188
rect -46 -281 -39 -274
rect -57 -293 -50 -286
rect -35 -363 -28 -356
rect -46 -375 -39 -368
rect -57 -387 -50 -380
rect 75 -139 82 -132
rect 35 -173 42 -166
rect 48 -183 55 -176
rect 11 -195 18 -188
rect 156 -53 163 -46
rect 167 -139 174 -132
rect 167 -171 174 -164
rect 156 -183 163 -176
rect 73 -195 80 -188
rect 145 -195 152 -188
rect 77 -233 84 -226
rect 35 -281 42 -274
rect 11 -293 18 -286
rect 89 -293 96 -286
rect 89 -326 96 -319
rect 48 -365 55 -358
rect 35 -375 42 -368
rect 11 -387 18 -380
rect 101 -422 108 -415
rect 77 -454 84 -447
rect 89 -465 96 -458
rect 101 -481 108 -474
rect 167 -293 174 -286
<< metal2 >>
rect -50 37 25 42
rect 82 33 145 38
rect -39 -49 25 -44
rect 82 -53 156 -48
rect -17 -135 25 -130
rect 82 -139 167 -134
rect 42 -171 167 -166
rect 55 -183 156 -178
rect -28 -195 11 -190
rect 80 -195 145 -190
rect -39 -281 35 -276
rect -50 -293 11 -288
rect -28 -363 48 -358
rect -39 -375 35 -370
rect -50 -387 11 -382
rect 79 -447 84 -233
rect 96 -293 167 -288
rect 91 -458 96 -326
rect 103 -474 108 -422
use 1INV  1INV_0
timestamp 1493152604
transform 1 0 49 0 1 20
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493152604
transform 1 0 49 0 1 -66
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493152604
transform 1 0 49 0 1 -152
box -49 -20 79 66
use 4NAND  4NAND_0
timestamp 1493152043
transform 1 0 18 0 1 -215
box -18 -55 110 43
use 3NAND  3NAND_0
timestamp 1493160834
transform 1 0 18 0 1 -313
box -18 -51 110 43
use 3NAND  3NAND_1
timestamp 1493160834
transform 1 0 18 0 1 -407
box -18 -51 110 43
use 3NAND  3NAND_2
timestamp 1493160834
transform 1 0 18 0 1 -501
box -18 -51 110 43
<< labels >>
rlabel metal1 -57 -552 -53 37 3 A
rlabel space -47 -553 -42 86 1 B
rlabel metal1 -35 -552 -31 86 1 C
rlabel space -24 -553 -20 86 1 D
<< end >>
