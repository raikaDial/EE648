magic
tech tsmc
timestamp 1493249588
<< metal1 >>
rect 0 86 4 92
rect 124 86 128 92
rect -57 44 -53 86
rect -57 -544 -53 37
rect -46 -42 -42 86
rect -46 -372 -42 -49
rect -35 -128 -31 86
rect -46 -544 -42 -379
rect -35 -544 -31 -135
rect -24 -188 -20 86
rect 32 37 36 41
rect 148 40 152 86
rect 71 33 75 37
rect 32 -49 36 -45
rect 66 -53 75 -49
rect 32 -135 36 -131
rect 66 -139 75 -135
rect 148 -188 152 33
rect 159 -46 163 86
rect 18 -195 25 -191
rect 42 -195 47 -191
rect -24 -278 -20 -195
rect 43 -225 62 -221
rect 37 -273 74 -269
rect 37 -277 41 -273
rect 18 -285 23 -281
rect 56 -285 74 -281
rect -24 -544 -20 -285
rect 60 -317 76 -313
rect 37 -367 86 -363
rect 18 -379 23 -375
rect 37 -376 41 -367
rect 148 -372 152 -195
rect 159 -278 163 -53
rect 170 -132 174 86
rect 170 -266 174 -139
rect 56 -379 86 -375
rect 60 -411 88 -407
rect 24 -443 62 -439
rect 24 -468 28 -443
rect 37 -454 74 -450
rect 37 -469 41 -454
rect 49 -473 86 -469
rect 56 -507 64 -503
rect 148 -544 152 -379
rect 159 -544 163 -285
rect 170 -360 174 -273
rect 170 -544 174 -367
<< m2contact >>
rect -57 37 -50 44
rect -46 -49 -39 -42
rect -35 -135 -28 -128
rect -46 -379 -39 -372
rect 25 37 32 44
rect 75 33 82 40
rect 145 33 152 40
rect 25 -49 32 -42
rect 75 -53 82 -46
rect 25 -135 32 -128
rect 75 -139 82 -132
rect 156 -53 163 -46
rect -24 -195 -17 -188
rect 11 -195 18 -188
rect 47 -195 54 -188
rect 145 -195 152 -188
rect 62 -228 69 -221
rect 74 -273 81 -266
rect -24 -285 -17 -278
rect 11 -285 18 -278
rect 74 -285 81 -278
rect 76 -320 83 -313
rect 86 -367 93 -360
rect 11 -379 18 -372
rect 167 -139 174 -132
rect 167 -273 174 -266
rect 156 -285 163 -278
rect 86 -379 93 -372
rect 145 -379 152 -372
rect 88 -411 95 -404
rect 62 -446 69 -439
rect 74 -454 81 -447
rect 86 -473 93 -466
rect 64 -507 71 -500
rect 167 -367 174 -360
<< metal2 >>
rect -50 37 25 42
rect 82 33 145 38
rect -39 -49 25 -44
rect 82 -53 156 -48
rect -28 -135 25 -130
rect 82 -139 167 -134
rect -17 -195 11 -190
rect 54 -195 145 -190
rect -17 -285 11 -280
rect -39 -379 11 -374
rect 64 -439 69 -228
rect 81 -273 167 -268
rect 81 -285 156 -280
rect 76 -447 81 -320
rect 93 -367 167 -362
rect 93 -379 145 -374
rect 88 -466 93 -411
rect 66 -551 71 -507
use 1INV  1INV_0
timestamp 1493248008
transform 1 0 49 0 1 20
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493248008
transform 1 0 49 0 1 -66
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493248008
transform 1 0 49 0 1 -152
box -49 -20 79 66
use 2NAND  2NAND_0
timestamp 1493246188
transform 1 0 16 0 1 -215
box -16 -47 112 43
use 3NAND  3NAND_0
timestamp 1493246171
transform 1 0 18 0 1 -305
box -18 -51 110 43
use 3NAND  3NAND_1
timestamp 1493246171
transform 1 0 18 0 1 -399
box -18 -51 110 43
use 3NAND  3NAND_2
timestamp 1493246171
transform 1 0 18 0 1 -493
box -18 -51 110 43
<< labels >>
rlabel metal1 -57 -544 -53 86 3 A
rlabel metal1 -46 -544 -42 86 1 B
rlabel metal1 -35 -544 -31 86 1 C
rlabel metal1 -24 -544 -20 86 1 D
rlabel metal1 0 86 4 92 5 Vdd
rlabel metal1 124 86 128 92 5 Gnd
rlabel metal2 66 -551 71 -546 1 Y
<< end >>
