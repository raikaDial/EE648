SEGMENT_C
* SPICE3 file created from seg_c.ext - technology: tsmc

.option scale=0.06u
.include mosistsmc180.sp

V_paprika_0 D Gnd PULSE(3.3 0 0 1n 1n 18n 40n)
V_paprika_1 C Gnd PULSE(3.3 0 0 1n 1n 38n 80n)
V_paprika_2 B Gnd PULSE(3.3 0 0 1n 1n 78n 160n)
V_paprika_3 A Gnd PULSE(3.3 0 0 1n 1n 158n 320n)
V_paprika_4 Vdd Gnd DC 3.3

M1000 Y m1_24_n475 Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=920 ps=422 
M1001 Vdd m1_37_n478 Y Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 Y m1_49_n481 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1003 x0/a_9_n26 m1_24_n475 Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=632 ps=286 
M1004 x0/a_22_n26 m1_37_n478 x0/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1005 Y m1_49_n481 x0/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1006 m1_49_n481 A Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1007 Vdd B m1_49_n481 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1008 m1_49_n481 C Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1009 x1/a_9_n26 A Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1010 x1/a_22_n26 B x1/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1011 m1_49_n481 C x1/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1012 m1_37_n478 A Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1013 Vdd B m1_37_n478 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1014 m1_37_n478 m1_35_n187 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1015 x2/a_9_n26 A Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1016 x2/a_22_n26 B x2/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1017 m1_37_n478 m1_35_n187 x2/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1018 m1_24_n475 C Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=0 ps=0 
M1019 Vdd m1_35_n187 m1_24_n475 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1020 m1_24_n475 m1_48_n190 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1021 Vdd m1_66_n195 m1_24_n475 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1022 x3/a_9_n30 C Gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1023 x3/a_22_n30 m1_35_n187 x3/a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1024 x3/a_35_n30 m1_48_n190 x3/a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1025 m1_24_n475 m1_66_n195 x3/a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1026 m1_35_n187 D Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1027 m1_35_n187 D Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1028 m1_48_n190 B Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1029 m1_48_n190 B Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1030 m1_66_n195 A Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1031 m1_66_n195 A Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
C0 m1_35_n187 m1_48_n190 4.8fF
C1 m1_37_n478 Y 0.0fF
C2 m1_49_n481 Y 0.0fF
C3 m1_24_n475 Vdd 0.8fF
C4 m1_37_n478 m1_49_n481 0.5fF
C5 m1_35_n187 Gnd 0.1fF
C6 m1_35_n187 m1_66_n195 0.0fF
C7 Gnd Y 0.1fF
C8 m1_37_n478 Gnd 0.1fF
C9 Gnd m1_49_n481 0.1fF
C10 Gnd m1_48_n190 0.1fF
C11 m1_66_n195 m1_48_n190 4.5fF
C12 m1_35_n187 m1_24_n475 0.1fF
C13 Gnd m1_66_n195 0.1fF
C14 m1_37_n478 m1_24_n475 1.4fF
C15 m1_24_n475 m1_49_n481 0.0fF
C16 m1_24_n475 m1_48_n190 0.0fF
C17 m1_35_n187 Vdd 0.3fF
C18 Gnd m1_24_n475 0.1fF
C19 Y Vdd 0.4fF
C20 m1_37_n478 Vdd 0.6fF
C21 m1_66_n195 m1_24_n475 0.0fF
C22 m1_49_n481 Vdd 0.5fF
C23 Vdd m1_48_n190 0.3fF
C24 m1_66_n195 Vdd 0.3fF
C25 m1_35_n187 m1_37_n478 0.0fF
C26 m1_66_n195 Gnd 1.6fF
C27 m1_48_n190 Gnd 1.6fF
C28 m1_35_n187 Gnd 2.2fF
C29 m1_24_n475 Gnd 0.3fF
C30 m1_37_n478 Gnd 0.4fF
C31 m1_49_n481 Gnd 0.5fF
C32 Gnd Gnd 2.6fF
C33 Y Gnd 0.1fF
C34 Vdd Gnd 6.1fF

** hspice subcircuit dictionary
* x0	3NAND_2
* x1	3NAND_1
* x2	3NAND_0
* x3	4NAND_0

.tran 1n 320n

.control
set filetype=ascii
run
write segC.txt A B C D Y
.endc
.end
