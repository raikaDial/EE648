* HSPICE file created from seg_c.ext - technology: tsmc

.option scale=0.06u

M1000 Y m1_24_n475 Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=920 ps=422 
M1001 Vdd m1_37_n478 Y Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 Y m1_49_n481 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1003 x0/a_9_n26 m1_24_n475 Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=632 ps=286 
M1004 x0/a_22_n26 m1_37_n478 x0/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1005 Y m1_49_n481 x0/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1006 m1_49_n481 A Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1007 Vdd m1_n46_n552 m1_49_n481 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1008 m1_49_n481 C Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1009 x1/a_9_n26 A Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1010 x1/a_22_n26 m1_n46_n552 x1/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1011 m1_49_n481 C x1/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1012 m1_37_n478 A Vdd Vdd pfet w=8 l=3
+ ad=152 pd=70 as=0 ps=0 
M1013 Vdd m1_n46_n552 m1_37_n478 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1014 m1_37_n478 m1_35_n187 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1015 x2/a_9_n26 A Gnd Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1016 x2/a_22_n26 m1_n46_n552 x2/a_9_n26 Gnd nfet w=12 l=3
+ ad=120 pd=44 as=0 ps=0 
M1017 m1_37_n478 m1_35_n187 x2/a_22_n26 Gnd nfet w=12 l=3
+ ad=108 pd=42 as=0 ps=0 
M1018 m1_24_n475 C Vdd Vdd pfet w=8 l=3
+ ad=160 pd=72 as=0 ps=0 
M1019 Vdd m1_35_n187 m1_24_n475 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1020 m1_24_n475 m1_48_n190 Vdd Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1021 Vdd m1_66_n195 m1_24_n475 Vdd pfet w=8 l=3
+ ad=0 pd=0 as=0 ps=0 
M1022 x3/a_9_n30 C Gnd Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1023 x3/a_22_n30 m1_35_n187 x3/a_9_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1024 x3/a_35_n30 m1_48_n190 x3/a_22_n30 Gnd nfet w=16 l=3
+ ad=160 pd=52 as=0 ps=0 
M1025 m1_24_n475 m1_66_n195 x3/a_35_n30 Gnd nfet w=16 l=3
+ ad=120 pd=50 as=0 ps=0 
M1026 m1_35_n187 m1_n24_n552 Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1027 m1_35_n187 m1_n24_n552 Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1028 m1_48_n190 m1_n46_n552 Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1029 m1_48_n190 m1_n46_n552 Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
M1030 m1_66_n195 A Vdd Vdd pfet w=8 l=3
+ ad=80 pd=36 as=0 ps=0 
M1031 m1_66_n195 A Gnd Gnd nfet w=4 l=3
+ ad=72 pd=36 as=0 ps=0 
C0 Vdd m1_n46_n552 0.5fF
C1 Gnd m1_24_n475 0.1fF
C2 Vdd m1_24_n475 0.8fF
C3 Vdd m1_n24_n552 0.1fF
C4 m1_66_n195 m1_48_n190 4.5fF
C5 m1_35_n187 m1_48_n190 4.8fF
C6 Gnd m1_37_n478 0.1fF
C7 Vdd m1_37_n478 0.6fF
C8 m1_48_n190 m1_24_n475 0.0fF
C9 m1_49_n481 m1_n46_n552 0.0fF
C10 Y m1_37_n478 0.0fF
C11 m1_49_n481 m1_24_n475 0.0fF
C12 Gnd Y 0.1fF
C13 Y Vdd 0.4fF
C14 Gnd m1_48_n190 0.1fF
C15 Vdd m1_48_n190 0.3fF
C16 m1_49_n481 m1_37_n478 0.5fF
C17 m1_66_n195 m1_35_n187 0.0fF
C18 m1_49_n481 Gnd 0.1fF
C19 m1_49_n481 Vdd 0.5fF
C20 m1_66_n195 m1_24_n475 0.0fF
C21 m1_49_n481 Y 0.0fF
C22 m1_n46_n552 m1_35_n187 0.1fF
C23 m1_35_n187 m1_24_n475 0.1fF
C24 m1_n24_n552 m1_n46_n552 0.0fF
C25 Gnd m1_66_n195 0.1fF
C26 Vdd m1_66_n195 0.3fF
C27 m1_35_n187 m1_37_n478 0.0fF
C28 Gnd m1_35_n187 0.1fF
C29 m1_n46_n552 m1_37_n478 0.0fF
C30 Vdd m1_35_n187 0.3fF
C31 m1_37_n478 m1_24_n475 1.4fF
C32 m1_66_n195 gnd! 1.6fF
C33 m1_48_n190 gnd! 1.6fF
C34 m1_n46_n552 gnd! 11.5fF
C35 m1_35_n187 gnd! 2.1fF
C36 m1_n24_n552 gnd! 5.3fF
C37 m1_24_n475 gnd! 0.3fF
C38 m1_37_n478 gnd! 0.4fF
C39 m1_49_n481 gnd! 0.5fF
C40 Gnd gnd! 2.6fF
C41 Y gnd! 0.1fF
C42 Vdd gnd! 5.5fF

** hspice subcircuit dictionary
* x0	3NAND_2
* x1	3NAND_1
* x2	3NAND_0
* x3	4NAND_0
