magic
tech tsmc
timestamp 1492555172
<< nwell >>
rect -13 17 30 50
<< ntransistor >>
rect 9 7 12 11
<< ptransistor >>
rect 9 25 12 33
<< ndiffusion >>
rect 7 7 9 11
rect 12 7 14 11
<< pdiffusion >>
rect 7 25 9 33
rect 12 25 14 33
<< ndcontact >>
rect -1 3 7 11
rect 14 3 22 11
<< pdcontact >>
rect -1 25 7 33
rect 14 25 22 33
<< nsubstratencontact >>
rect 14 40 22 48
<< polysilicon >>
rect 9 33 12 37
rect 9 20 12 25
rect -5 17 12 20
rect 9 11 12 17
rect 9 3 12 7
<< polycontact >>
rect -13 17 -5 25
<< metal1 >>
rect -47 58 -43 66
rect -47 54 20 58
rect -47 -20 -43 54
rect 16 48 20 54
rect -1 40 14 46
rect -1 33 4 40
rect 17 11 22 25
rect 1 -2 5 3
rect 71 -2 75 66
rect 1 -6 75 -2
rect 71 -20 75 -6
<< labels >>
rlabel metal1 -47 -14 -43 66 3 Vdd
rlabel metal1 71 -14 75 66 7 Gnd
rlabel polycontact -13 17 -5 25 1 A
rlabel metal1 17 11 22 25 1 Y
<< end >>
