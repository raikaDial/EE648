magic
tech tsmc
timestamp 1493253861
<< metal1 >>
rect -57 -213 -53 86
rect -46 -128 -42 86
rect -35 -42 -31 86
rect -24 44 -20 86
rect 32 37 39 41
rect -57 -454 -53 -220
rect -46 -344 -42 -135
rect -57 -490 -53 -461
rect -46 -466 -42 -351
rect -35 -356 -31 -49
rect -46 -491 -42 -473
rect -35 -490 -31 -363
rect -24 -368 -20 37
rect 69 36 75 40
rect 29 -49 36 -45
rect 69 -50 75 -46
rect 32 -135 40 -131
rect 70 -137 75 -132
rect 32 -219 40 -215
rect 148 -217 152 86
rect 159 -130 163 86
rect 170 -43 174 86
rect 181 43 185 86
rect 70 -224 75 -219
rect 24 -277 28 -259
rect 37 -275 42 -269
rect 54 -278 78 -275
rect 148 -278 152 -224
rect 159 -262 163 -137
rect 170 -250 174 -50
rect 54 -279 72 -278
rect 59 -314 76 -309
rect 36 -368 41 -363
rect 50 -367 54 -353
rect 148 -367 152 -285
rect 18 -374 25 -370
rect 69 -374 88 -369
rect -24 -491 -20 -375
rect 73 -409 88 -408
rect 72 -412 88 -409
rect 72 -414 73 -412
rect 0 -465 4 -448
rect 50 -460 100 -455
rect 37 -465 41 -461
rect 50 -466 55 -460
rect 18 -472 25 -468
rect 69 -473 100 -467
rect 148 -490 152 -374
rect 159 -491 163 -269
rect 170 -466 174 -257
rect 181 -454 185 36
rect 170 -490 174 -473
rect 181 -491 185 -461
rect 73 -511 100 -506
rect 23 -548 100 -542
rect 23 -563 29 -548
rect 37 -558 88 -554
rect 37 -565 41 -558
rect 54 -571 76 -566
<< m2contact >>
rect -24 37 -17 44
rect 25 37 32 44
rect -35 -49 -28 -42
rect -46 -135 -39 -128
rect -57 -220 -50 -213
rect -46 -351 -39 -344
rect -57 -461 -50 -454
rect -35 -363 -28 -356
rect -46 -473 -39 -466
rect 75 36 82 43
rect 22 -49 29 -42
rect 75 -50 82 -43
rect 25 -135 32 -128
rect 75 -137 82 -130
rect 25 -220 32 -213
rect 178 36 185 43
rect 168 -50 175 -43
rect 156 -137 163 -130
rect 75 -224 82 -217
rect 145 -224 152 -217
rect 23 -259 30 -252
rect 36 -269 43 -262
rect 167 -257 174 -250
rect 156 -269 163 -262
rect 72 -285 79 -278
rect 145 -285 152 -278
rect 76 -314 83 -307
rect 48 -353 55 -346
rect 35 -363 42 -356
rect -24 -375 -17 -368
rect 11 -375 18 -368
rect 88 -374 95 -367
rect 146 -374 153 -367
rect 88 -412 95 -405
rect 36 -461 43 -454
rect 100 -461 107 -454
rect 11 -473 18 -466
rect 100 -473 107 -466
rect 178 -461 185 -454
rect 168 -473 175 -466
rect 100 -512 107 -505
rect 100 -548 107 -541
rect 88 -559 95 -552
rect 76 -571 83 -564
<< metal2 >>
rect -17 37 25 42
rect 82 36 178 41
rect -28 -49 22 -44
rect 82 -50 168 -44
rect -39 -135 25 -130
rect 82 -137 156 -132
rect -50 -219 25 -214
rect 82 -224 145 -219
rect 30 -257 167 -252
rect 43 -269 156 -263
rect 79 -285 145 -279
rect -39 -351 48 -346
rect -28 -363 35 -358
rect -17 -375 11 -370
rect -50 -461 36 -456
rect -39 -473 11 -468
rect 78 -564 83 -314
rect 95 -374 146 -369
rect 90 -552 95 -412
rect 107 -461 178 -456
rect 107 -473 168 -468
rect 101 -541 106 -512
use 1INV  1INV_0
timestamp 1493152604
transform 1 0 49 0 1 20
box -49 -20 79 66
use 1INV  1INV_1
timestamp 1493152604
transform 1 0 49 0 1 -66
box -49 -20 79 66
use 1INV  1INV_2
timestamp 1493152604
transform 1 0 49 0 1 -152
box -49 -20 79 66
use 1INV  1INV_3
timestamp 1493152604
transform 1 0 49 0 1 -238
box -49 -20 79 66
use 3NAND  3NAND_0
timestamp 1492655848
transform 1 0 18 0 1 -301
box -18 -51 110 43
use 4NAND  4NAND_0
timestamp 1493152043
transform 1 0 18 0 1 -395
box -18 -55 110 43
use 4NAND  4NAND_1
timestamp 1493152043
transform 1 0 18 0 1 -493
box -18 -55 110 43
use 3NAND  3NAND_1
timestamp 1492655848
transform 1 0 18 0 1 -591
box -18 -51 110 43
<< end >>
